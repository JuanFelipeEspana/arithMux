`timescale 1 ns/ 10 ps
module fullAdder4b_tb();
   reg[3:0] a_tb, b_tb;
   wire[3:0] sum_tb;
   wire      cout_tb;

   fullAdder4b DUT (.a(a_tb),.b(b_tb),.cin(1'b0),.sum(sum_tb),.cout(cout_tb));

   initial
     begin
	a_tb = 4'b0000;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0001;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0010;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0011;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0100;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0101;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0110;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b0111;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1000;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1001;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1010;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1011;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1100;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1101;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1110;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	a_tb = 4'b1111;
	b_tb = 4'b0000;
	# 200;
	b_tb = 4'b0001;
	# 200;
	b_tb = 4'b0010;
	# 200;
	b_tb = 4'b0011;
	# 200;
	b_tb = 4'b0100;
	# 200;
	b_tb = 4'b0101;
	# 200;
	b_tb = 4'b0110;
	# 200;
	b_tb = 4'b0111;
	# 200;
	b_tb = 4'b1000;
	# 200;
	b_tb = 4'b1001;
	# 200;
	b_tb = 4'b1010;
	# 200;
	b_tb = 4'b1011;
	# 200;
	b_tb = 4'b1100;
	# 200;
	b_tb = 4'b1101;
	# 200;
	b_tb = 4'b1110;
	# 200;
	b_tb = 4'b1111;
	# 200;
	$stop;
     end // initial begin
endmodule
   
